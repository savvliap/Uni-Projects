library verilog;
use verilog.vl_types.all;
entity counter4bit_tb is
end counter4bit_tb;
